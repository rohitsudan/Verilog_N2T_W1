`timescale 1ns/10ps
module testbench_simple;
parameter width = 16;
reg [width-1:0] in0,in1,in2,in3,in4,in5,in6,in7;
reg [2:0] sel;
wire [width-1:0] out;
mux8to1_16bit mymux(in0,in1,in2,in3,in4,in5,in6,in7,sel,out);
initial
begin
	$dumpfile("testbench_simple.vcd");//the name of the .vcd file should be as the same as the testbecnh file
	$dumpvars(0,testbench_simple);
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b000;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b001;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b010;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b011;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b100;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b101;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b110;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b111;
	#1;
	in0='b1111111111111111;
	in1='b0000000000000000;
	in2='b1111111000000000;
	in3='b0000000111111111;
	in4='b0001000111111111;
	in5='b0000000111110111;
	in6='b0100000111110111;
	in7='b1100000111111111;
	sel='b111;
        $finish;
end
endmodule

module orgate(in0,in1,out);
input in0,in1;
output out;
//and and1(out,in0,in1);
assign out = in0 | in1; // please check out under what this comes

endmodule
